typedef uvm_sequencer#(wr_tx) wr_sqr;

typedef uvm_sequencer#(rd_tx) rd_sqr;


// class wr_sqr extends uvm_sequencer #(wr_tx);
  
//   `uvm_component_utils(wr_sqr)
  
//   function new(string name = "", uvm_component parent = null);
//     super.new(name, parent);
//   endfunction
  
//   function void build_phase (uvm_phase phase);
//     super.build_phase(phase);
    
//   endfunction
  
// endclass